module play