module play 

import primitives

fn test_player() {
	base := init_basic_stats(primitives.phys(2))
	println(base)
	atts := base.init_attributes()
	println(atts)
}