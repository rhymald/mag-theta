module play 

// import primitives

fn test_player() {
	base := init_basic_stats()
	println(base)
	atts := base.init_attributes()
	println(atts)
}