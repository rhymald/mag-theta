module funcs

import time