module play

import funcs

struct Attributes {
	toughness f64
	vitality f64
	stamina f64
	power f64
}

fn (base BasicStats) init_attributes() Attributes {
	return Attributes{
		toughness: funcs.round((1 + base.body.c + 2*base.body.d + base.body.a) / 3)
		power: funcs.round((1 + base.body.a + 2*base.body.d + base.body.c) / 3)
		vitality: funcs.round(100 + (1 + base.body.a + 2*base.body.c ) / 3)
		stamina: funcs.round(100 + (1 + 2*base.body.c + base.body.d) / 3)
	}
}