module funcs

fn test_me() {
	for _ in 0..12 {
		print(round(init_f64()))
		print(' ')
	}
}