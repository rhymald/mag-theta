module funcs